library verilog;
use verilog.vl_types.all;
entity eightBusInterface_tb is
end eightBusInterface_tb;
