library verilog;
use verilog.vl_types.all;
entity tb_inputWrapper is
end tb_inputWrapper;
