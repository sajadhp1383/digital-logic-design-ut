library verilog;
use verilog.vl_types.all;
entity tb_outputWrapper is
end tb_outputWrapper;
