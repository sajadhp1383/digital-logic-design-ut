`timescale 1ns/1ns

module myNOT(input a,output w);
	supply1 vdd;
	supply0 gnd;
	pmos #(4,7,9) T1(w,vdd,a);
	nmos #(3,5,7) T2(w,gnd,a);
endmodule;
